module S011HD1P_X256Y2D32(
    Q, CLK, CEN, WEN, A, D
);
parameter Bits = 32;
parameter Word_Depth = 512;
parameter Add_Width = 9;
parameter Wen_Width = 32;

output reg [Bits-1:0] Q;
input                 CLK;
input                 CEN;
input                 WEN;
input [Add_Width-1:0] A;
input [Bits-1:0]      D;

wire cen  = ~CEN;
wire wen  = ~WEN;

reg [Bits-1:0] ram [0:Word_Depth-1];
always @(posedge CLK) begin
    if(cen && wen) begin
        ram[A] <= D;
    end
    Q <= cen && !wen ? ram[A] : {4{$random}};
end

endmodule