// combine mapping and vga_ctrl_axi

module vga_ctrl(
    input clock,
	input resetn,
    input         io_master_awready,
    output        io_master_awvalid,
    output [31:0] io_master_awaddr,
    output [3:0]  io_master_awid,
    output [7:0]  io_master_awlen,
    output [2:0]  io_master_awsize,
    output [1:0]  io_master_awburst,
    input         io_master_wready,
    output        io_master_wvalid,
    output [63:0] io_master_wdata,
    output [7:0]  io_master_wstrb,
    output        io_master_wlast,
    output        io_master_bready,
    input         io_master_bvalid,
    input  [1:0]  io_master_bresp,
    input  [3:0]  io_master_bid,
    input         io_master_arready,
    output        io_master_arvalid,
    output [31:0] io_master_araddr,
    output [3:0]  io_master_arid,
    output [7:0]  io_master_arlen,
    output [2:0]  io_master_arsize,
    output [1:0]  io_master_arburst,
    output        io_master_rready,
    input         io_master_rvalid,
    input  [1:0]  io_master_rresp,
    input  [63:0] io_master_rdata,
    input         io_master_rlast,
    input  [3:0]  io_master_rid,

    output        io_slave_map_awready,
    input         io_slave_map_awvalid,
    input  [31:0] io_slave_map_awaddr,
    input  [3:0]  io_slave_map_awid,
    input  [7:0]  io_slave_map_awlen,
    input  [2:0]  io_slave_map_awsize,
    input  [1:0]  io_slave_map_awburst,
    output        io_slave_map_wready,
    input         io_slave_map_wvalid,
    input  [63:0] io_slave_map_wdata,
    input  [7:0]  io_slave_map_wstrb,
    input         io_slave_map_wlast,
    input         io_slave_map_bready,
    output        io_slave_map_bvalid,
    output [1:0]  io_slave_map_bresp,
    output [3:0]  io_slave_map_bid,
    output        io_slave_map_arready,
    input         io_slave_map_arvalid,
    input  [31:0] io_slave_map_araddr,
    input  [3:0]  io_slave_map_arid,
    input  [7:0]  io_slave_map_arlen,
    input  [2:0]  io_slave_map_arsize,
    input  [1:0]  io_slave_map_arburst,
    input         io_slave_map_rready,
    output        io_slave_map_rvalid,
    output [1:0]  io_slave_map_rresp,
    output [63:0] io_slave_map_rdata,
    output        io_slave_map_rlast,
    output [3:0]  io_slave_map_rid,

    output        io_slave_vga_awready,
    input         io_slave_vga_awvalid,
    input  [31:0] io_slave_vga_awaddr,
    input  [3:0]  io_slave_vga_awid,
    input  [7:0]  io_slave_vga_awlen,
    input  [2:0]  io_slave_vga_awsize,
    input  [1:0]  io_slave_vga_awburst,
    output        io_slave_vga_wready,
    input         io_slave_vga_wvalid,
    input  [63:0] io_slave_vga_wdata,
    input  [7:0]  io_slave_vga_wstrb,
    input         io_slave_vga_wlast,
    input         io_slave_vga_bready,
    output        io_slave_vga_bvalid,
    output [1:0]  io_slave_vga_bresp,
    output [3:0]  io_slave_vga_bid,
    output        io_slave_vga_arready,
    input         io_slave_vga_arvalid,
    input  [31:0] io_slave_vga_araddr,
    input  [3:0]  io_slave_vga_arid,
    input  [7:0]  io_slave_vga_arlen,
    input  [2:0]  io_slave_vga_arsize,
    input  [1:0]  io_slave_vga_arburst,
    input         io_slave_vga_rready,
    output        io_slave_vga_rvalid,
    output [1:0]  io_slave_vga_rresp,
    output [63:0] io_slave_vga_rdata,
    output        io_slave_vga_rlast,
    output [3:0]  io_slave_vga_rid,

    output hsync,
	output vsync,
	output [3:0]vga_r,
	output [3:0]vga_g,
	output [3:0]vga_b

);

    wire [31:0] offset;

    vga_ctrl_comb vga(
        .clock(clock),
        .resetn(resetn),
        .io_master_awready(1'b0),
        // .io_master_awvalid,
        // .io_master_awaddr,
        // .io_master_awid,
        // .io_master_awlen,
        // .io_master_awsize,
        // .io_master_awburst,
        .io_master_wready(1'b0),
        // .io_master_wvalid,
        // .io_master_wdata,
        // .io_master_wstrb,
        // .io_master_wlast,
        .io_master_bready(1'b0),
        // .io_master_bvalid,
        // .io_master_bresp,
        // .io_master_bid,
        .io_master_arready(io_master_arready),
        .io_master_arvalid(io_master_arvalid),
        .io_master_araddr(io_master_araddr),
        .io_master_arid(io_master_arid),
        .io_master_arlen(io_master_arlen),
        .io_master_arsize(io_master_arsize),
        .io_master_arburst(io_master_arburst),
        .io_master_rready(io_master_rready),
        .io_master_rvalid(io_master_rvalid),
        .io_master_rresp(io_master_rresp),
        .io_master_rdata(io_master_rdata),
        .io_master_rlast(io_master_rlast),
        .io_master_rid(io_master_rid),

        .io_slave_awready(io_slave_vga_awready),
        .io_slave_awvalid(io_slave_vga_awvalid),
        .io_slave_awaddr(io_slave_vga_awaddr),
        .io_slave_awid(io_slave_vga_awid),
        .io_slave_awlen(io_slave_vga_awlen),
        .io_slave_awsize(io_slave_vga_awsize),
        .io_slave_awburst(io_slave_vga_awburst),
        .io_slave_wready(io_slave_vga_wready),
        .io_slave_wvalid(io_slave_vga_wvalid),
        .io_slave_wdata(io_slave_vga_wdata),
        .io_slave_wstrb(io_slave_vga_wstrb),
        .io_slave_wlast(io_slave_vga_wlast),
        .io_slave_bready(io_slave_vga_bready),
        .io_slave_bvalid(io_slave_vga_bvalid),
        .io_slave_bresp(io_slave_vga_bresp),
        .io_slave_bid(io_slave_vga_bid),
        .io_slave_arready(io_slave_vga_arready),
        .io_slave_arvalid(io_slave_vga_arvalid),
        .io_slave_araddr(io_slave_vga_araddr),
        .io_slave_arid(io_slave_vga_arid),
        .io_slave_arlen(io_slave_vga_arlen),
        .io_slave_arsize(io_slave_vga_arsize),
        .io_slave_arburst(io_slave_vga_arburst),
        .io_slave_rready(io_slave_vga_rready),
        .io_slave_rvalid(io_slave_vga_rvalid),
        .io_slave_rresp(io_slave_vga_rresp),
        .io_slave_rdata(io_slave_vga_rdata),
        .io_slave_rlast(io_slave_vga_rlast),
        .io_slave_rid(io_slave_vga_rid),

        .io_offset(offset),
        .hsync(hsync),
        .vsync(vsync),
        .vga_r(vga_r),
        .vga_g(vga_g),
        .vga_b(vga_b)
    );

    Mapping map(
        .clock(clock),
        .reset(~resetn),
        .io_map_in_awready(io_slave_map_awready),
        .io_map_in_awvalid(io_slave_map_awvalid),
        .io_map_in_awaddr(io_slave_map_awaddr),
        .io_map_in_awid(io_slave_map_awid),
        .io_map_in_awlen(io_slave_map_awlen),
        .io_map_in_awsize(io_slave_map_awsize),
        .io_map_in_awburst(io_slave_map_awburst),
        .io_map_in_wready(io_slave_map_wready),
        .io_map_in_wvalid(io_slave_map_wvalid),
        .io_map_in_wdata(io_slave_map_wdata),
        .io_map_in_wstrb(io_slave_map_wstrb),
        .io_map_in_wlast(io_slave_map_wlast),
        .io_map_in_bready(io_slave_map_bready),
        .io_map_in_bvalid(io_slave_map_bvalid),
        .io_map_in_bresp(io_slave_map_bresp),
        .io_map_in_bid(io_slave_map_bid),
        .io_map_in_arready(io_slave_map_arready),
        .io_map_in_arvalid(io_slave_map_arvalid),
        .io_map_in_araddr(io_slave_map_araddr),
        .io_map_in_arid(io_slave_map_arid),
        .io_map_in_arlen(io_slave_map_arlen),
        .io_map_in_arsize(io_slave_map_arsize),
        .io_map_in_arburst(io_slave_map_arburst),
        .io_map_in_rready(io_slave_map_rready),
        .io_map_in_rvalid(io_slave_map_rvalid),
        .io_map_in_rresp(io_slave_map_rresp),
        .io_map_in_rdata(io_slave_map_rdata),
        .io_map_in_rlast(io_slave_map_rlast),
        .io_map_in_rid(io_slave_map_rid),
        .io_offset(offset),
        .io_map_out_awready(io_master_awready),
        .io_map_out_awvalid(io_master_awvalid),
        .io_map_out_awaddr(io_master_awaddr),
        .io_map_out_awid(io_master_awid),
        .io_map_out_awlen(io_master_awlen),
        .io_map_out_awsize(io_master_awsize),
        .io_map_out_awburst(io_master_awburst),
        .io_map_out_wready(io_master_wready),
        .io_map_out_wvalid(io_master_wvalid),
        .io_map_out_wdata(io_master_wdata),
        .io_map_out_wstrb(io_master_wstrb),
        .io_map_out_wlast(io_master_wlast),
        .io_map_out_bready(io_master_bready),
        .io_map_out_bvalid(io_master_bvalid),
        .io_map_out_bresp(io_master_bresp),
        .io_map_out_bid(io_master_bid),
        .io_map_out_arready(0),
        // .io_map_out_arvalid,
        // .io_map_out_araddr,
        // .io_map_out_arid,
        // .io_map_out_arlen,
        // .io_map_out_arsize,
        // .io_map_out_arburst,
        // .io_map_out_rready,
        .io_map_out_rvalid(1'b0),
        .io_map_out_rresp(2'b0),
        .io_map_out_rdata(32'b0),
        .io_map_out_rlast(1'b0),
        .io_map_out_rid(4'b0)
    );

endmodule

